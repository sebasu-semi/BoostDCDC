* Extracted by KLayout

.SUBCKT TOP SW Vg Vo GND
M$1 GND Vg SW GND NCHOR1EX L=2U W=400U AS=404P AD=404P PS=606U PD=606U
M$101 SW Vo Vo SW PCHOR1EX L=2U W=660U AS=666.6P AD=666.6P PS=868.6U PD=868.6U
.ENDS TOP
